library IEEE; use IEEE.STD_LOGIC_1164.all;

entity flopra is
    port(ck: in STD_LOGIC;
         reset: in STD_LOGIC;
         d: in STD_LOGIC_VECTOR(3 downto 0);
         q: out STD_LOGIC_VECTOR(3 downto 0));
end;

architecture asynchronous of flopra is
begin
    process(ck, reset) begin
        if reset = '1' then
            q <= "0000";
        elsif ck' event and ck = '1' then
            q <= d;
        end if;
    end process;
end;
